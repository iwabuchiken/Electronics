CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
330 240 30 200 9
40 112 1560 1118
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
31 C:\WORKS\PROGRAMS\CM60S\BOM.DAT
0 7
40 112 1560 1118
144179218 0
0
6 Title:
5 Name:
0
0
0
6
9 Resistor~
219 590 594 0 1 5
0 0
0
0 0 864 180
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8953 0 0
0
0
7 Ground~
168 657 629 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
7 AD8561~
219 644 457 0 1 17
0 0
0
0 0 2880 90
5 LM385
30 -4 65 4
2 U1
41 -14 55 -6
0
0
29 %D %1 %2 %3 %4 %5 %6 %7 %8 %S
0
0
4 DIP8
17

0 2 3 1 4 5 6 7 8 2
3 1 4 5 6 7 8 0
88 0 0 0 1 1 0 0
1 U
3618 0 0
0
0
11 NLI Source~
204 859 456 0 1 5
0 0
0
0 0 16576 0
5 100mA
13 0 48 8
5 NLIs2
13 -10 48 -2
0
0
13 %D %1 %2 I=%L
0
0
0
5

0 1 2 1 2 0
66 0 0 0 0 0 0 0
4 NLIs
6153 0 0
0
0
11 NLI Source~
204 455 446 0 1 5
0 0
0
0 0 16448 0
5 100mA
13 0 48 8
5 NLIs1
13 -10 48 -2
0
0
13 %D %1 %2 I=%L
0
0
0
5

0 1 2 1 2 0
66 0 0 0 0 0 0 0
4 NLIs
5394 0 0
0
0
12 NPN Trans:B~
219 610 378 0 1 7
0 0
0
0 0 832 0
3 NPN
17 0 38 8
2 Q1
21 -10 35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
7734 0 0
0
0
5
1 1 0 0 0 0 0 3 1 0 0 3
639 486
639 594
608 594
3 2 0 0 0 16 0 3 1 0 0 5
630 486
630 554
565 554
565 594
572 594
4 1 0 0 0 0 0 3 2 0 0 2
657 486
657 623
2 2 0 0 0 0 0 4 5 0 0 4
859 477
859 473
455 473
455 467
1 1 0 0 0 0 0 5 4 0 0 4
455 425
455 432
859 432
859 435
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
